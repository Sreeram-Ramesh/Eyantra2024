// Module: Ripple Carry Adder
// Inputs: A[0:1], B[0:1], Cin
// Outputs: Sum[0:1], Cout

module ripple_carry_adder(in_1, in_2, c_in, sum, c_out);

	input [1:0] in_1, in_2;
	input c_in;
	output [1:0] sum;
	output c_out;
	
	wire c1;
	
	full_adder fa1(
		
		.in_1(in_1[0]),
		.in_2(in_2[0]),
		.c_in(c_in),
		.sum(sum[0]),
		.c_out(c1)
	
	);
	
	full_adder fa2(
	
		.in_1(in_1[1]),
		.in_2(in_2[1]),
		.c_in(c1),
		.sum(sum[1]),
		.c_out(c_out)
	);

endmodule